module mac_core(
    input wire clk,
    input wire reset_n,
    input wire [15:0] data_in,
    input wire wr_en,
    input wire rd_en,
    output wire [15:0] output,
    output wire output_ready
);
endmodule