module clock_generator(
    input wire clk_in,
    output wire clk_out
);
endmodule