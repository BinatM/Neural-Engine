module test_generator(
    input wire clk,
    input wire reset_n,
    input wire start,
    input wire [15:0] test_data_in,
    output wire [15:0] data_out,
    output wire [10:0] address,
    output wire wr_en,
    output wire rd_en,
    output wire chip_sel
);
endmodule