module control_unit(
    input wire clk,
    input wire reset_n,
    input wire start,
    output wire wr_en,
    output wire rd_en,
    output wire output_ready
);
endmodule